module MetroFSM
// ???????? CODE_BITS ???????? ?????????? ??? ??? ???????? ????
// ???????? MONEY_BITS ???????? ?????????? ??? ??? ???????? ????? 
#(parameter CODE_BITS = 6, MONEY_BITS = 14)
// clk - ???????? ??????
// ena - ?????????? ?????
// res - ?????????? ?????
// reset - ??????????? ?????
// code - ??? ??? ????????
// indicators - ??????????
(input wire clk, ena, res, reset, input wire isCardAttached,
input wire [MONEY_BITS-1:0] currentBalance, input wire [CODE_BITS-1:0] code,
output reg permission,
output wire [6:0] indicators0, [6:0] indicators1, [6:0] indicators2, [6:0] indicators3);
// ?????????
parameter INITIAL_STATE = 0; 
parameter CARD_WAITING_STATE = 1; 
parameter CARD_READING_STATE = 2; 
parameter CARD_DISPLAY_STATE = 3; 
parameter ENTRY_PERMIT_STATE = 4;
parameter CARD_READING_ERROR_STATE = 5;
// ??????????
reg [3:0] in4 [3:0];
MetroCoder cdr1 (.in4(in4[0]), .out7(indicators0)); 
MetroCoder cdr2 (.in4(in4[1]), .out7(indicators1)); 
MetroCoder cdr3 (.in4(in4[2]), .out7(indicators2)); 
MetroCoder cdr4 (.in4(in4[3]), .out7(indicators3));
// ?????????, ????, ???. ?????????? ? ????????? ???????
reg [2:0] state = INITIAL_STATE; 
reg [3:0] cnt = 0;
reg s;
reg [CODE_BITS-2:0] i, endi = CODE_BITS >> 1;
reg [MONEY_BITS-1:0] price = 6'b101101, newBalance;
// ?????????? ??????????? ???????
always@ (posedge clk or negedge reset) 
	if (!reset) begin
		state <= INITIAL_STATE;
		cnt <= 4'd0;
	end
// ?????? ???? ?????????
always@ (posedge clk or posedge reset) 
	if (res) begin
		state <= INITIAL_STATE;
		cnt <= 4'd0;
	end
	else case (state)
		INITIAL_STATE: begin
		// ??????? ? ????????? ???????? 
		in4[0] = 4'b1010; //			'_' 
		in4[1] = 4'b1010; //		'_' 
		in4[2] = 4'b1010; //	'_' 
		in4[3] = 4'b1010; // '_' 
		permission = 1'b0;
		state <= CARD_WAITING_STATE;
	end
	CARD_WAITING_STATE:
		// ??????? ? ??????, ???? 2 ????? ?????? 
		if (cnt == 4'd2) begin
			in4[0] = 4'b1011; //			'?' 
			in4[1] = 4'b1011; //		'?' 
			in4[2] = 4'b1011; //	'?' 
			in4[3] = 4'b1011; // '?'
			state <= CARD_READING_STATE;
		end
	CARD_READING_STATE:
	// ???? ????? ?? ?????????, ?? ??????? ? ??????????? ?????? 
	if (!isCardAttached) begin
		in4[0] = 4'b1100; //			'E' 
		in4[1] = 4'b1100; //		'E' 
		in4[2] = 4'b1100; //	'E' 
		in4[3] = 4'b1100; //'E'
		state <= CARD_READING_ERROR_STATE;
	end
	// ??????? ? ????????, ???? 2 ????? ?????? 
	else if (cnt == 4'd4) begin
		// ???????? ???? ? ???????
		// ???????? ????: ??? ??????, ???? ??????? ???? ???? ?????????????? ??????? ?????
		// ?. ?. ???? ???? n, ..., n/2 ?????????????? n/2-1, ..., 0 
		s = 1;
		for (i = 0; i < endi; i = i + 1'b1)
		s = s & (code[i] ^ code[i + endi]);
		// ???????? ???????: ???? ??????, ?? ????? ? ???????
		if (currentBalance < price || !s) 
			begin in4[0] = 4'b1100; //			'E' 
			in4[1] = 4'b1100; //		'E' 
			in4[2] = 4'b1100; //	'E'
			in4[3] = 4'b1100; // 'E'
			state <= CARD_READING_ERROR_STATE;
		end
		else begin
		// ??????? ????? ?? ???????? ? ?????????? ??? ??????????? 
		newBalance = currentBalance - price;
		i = 0;
		while (newBalance >= 1000) begin 
			newBalance = newBalance - 1000; 
			i = i + 1;
		end
		in4[3] = i; 
		i = 0;
		while (newBalance >= 100) begin 
			newBalance = newBalance - 100; 
			i = i + 1;
		end
		in4[2] = i; 
		i = 0;
		while (newBalance >= 10) begin 
			newBalance = newBalance - 10; 
			i = i + 1;
		end
		in4[1] = i;
		in4[0] = newBalance;
		state <= CARD_DISPLAY_STATE;
		end
	end
CARD_DISPLAY_STATE:
	// ??????? ? ?????????? ?????, ???? 3 ????? ?????? 
	if (cnt == 4'd7) begin
		permission <= 1'b1;
		state <= ENTRY_PERMIT_STATE;
	end
	ENTRY_PERMIT_STATE: begin
		in4[0] = 4'b1010; //			'_' 
		in4[1] = 4'b1010; //		'_' 
		in4[2] = 4'b1010; //	'_' 
		in4[3] = 4'b1010; // '_' 
		permission = 1'b0;
		state <= CARD_WAITING_STATE;
	end
	CARD_READING_ERROR_STATE: begin 
		in4[0] = 4'b1010; //			'_' 
		in4[1] = 4'b1010; //		'_' 
		in4[2] = 4'b1010; //	'_' 
		in4[3] = 4'b1010; // '_'
		state <= CARD_WAITING_STATE;
	end
endcase
// ?????? ???????? ?????? ?????????
always@ (posedge clk) 
	if (res) begin
		state <= INITIAL_STATE;
		cnt <= 4'd0;
	end
	else if (ena) case (state)
		INITIAL_STATE: begin
			cnt <= 4'd0;
		end
	CARD_WAITING_STATE: begin
		cnt <= (isCardAttached ? cnt + 4'd1 : 4'd0);
	end
	CARD_READING_STATE: begin
		cnt <= cnt + 4'd1;
	end
	CARD_DISPLAY_STATE: begin
		cnt <= cnt + 4'd1;
	end
	ENTRY_PERMIT_STATE: begin
		cnt <= 4'd0;
	end
	CARD_READING_ERROR_STATE: begin
		cnt <= 4'd0;
	end
	endcase 
endmodule


